----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/05/2024 02:52:54 PM
-- Design Name: 
-- Module Name: D_FF_Sim - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity D_FF_Sim is
--  Port ( );
end D_FF_Sim;

architecture Behavioral of D_FF_Sim is

Component D_FF is
    Port ( D : in STD_LOGIC;
           Res : in STD_LOGIC;
           Clk : in STD_LOGIC;
           Q : out STD_LOGIC;
           Qbar : out STD_LOGIC);
end component;

SIGNAL d, res, clk : STD_LOGIC;
SIGNAL q, qbar :  STD_LOGIC;

begin

UUT: D_FF port map(
    D => d, 
    Res => res,
    Clk => clk,
    Q => q,
    Qbar => qbar);
    
process
begin
    
    clk <= '0';
    d <= '1';
    res <= '0';
    wait for 10ns;
    clk <= '1';
    
    wait for 40ns;
    clk <= '0';
    
    wait for 50ns;
    clk <= '1';
    d <= '0';
    
    wait for 100ns;
    
    clk <= '0';
    res <= '0';
    
    wait for 100ns;
        
    d <= '1';
    
    wait for 100ns;
            
    clk <= '1';
    res <= '0';
    
    wait for 100ns;
                
    clk <= '0';
    d <= '1';
    wait for 100ns;
                
    d <= '0';
    
    wait for 100ns;
                
    res <= '1';
    
    wait;
end process;

end Behavioral;
